package Environment;
  `include "command.sv"
  `include "driver.sv" 
  `include "result.sv"
  `include "monitor.sv"
  `include "environment.sv"
endpackage : Environment

